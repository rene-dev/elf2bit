library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library work;
use work.mpsoc_config.all;
use work.zpu_config.all;



entity dualport_ram is
	generic(addrBitBRAM		: integer := 1);
	port(clk				: in  std_logic;
		 memAWriteEnable	: in  std_logic;
		 memAAddr			: in  std_logic_vector(addrBitBRAM downto minAddrBit);		-- 13 downto 2
		 memAWrite			: in  std_logic_vector(wordSize - 1 downto 0);
		 memARead			: out std_logic_vector(wordSize - 1 downto 0);
		 memBWriteEnable	: in  std_logic;
		 memBAddr			: in  std_logic_vector(addrBitBRAM downto minAddrBit);
		 memBWrite			: in  std_logic_vector(wordSize - 1 downto 0);
		 memBRead			: out std_logic_vector(wordSize - 1 downto 0));
end dualport_ram;



architecture behave_dualport_ram1 of dualport_ram is

begin

	RAMB16_S18_S18_inst1: RAMB16_S18_S18
		generic map (
INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000")
		port map (DOA => memARead(31 downto 16),
				  DOB => memBRead(31 downto 16),
				  DOPA => open,
				  DOPB => open,
				  ADDRA => memAAddr(addrBitBRAM downto minAddrBit),
				  ADDRB => memBAddr(addrBitBRAM downto minAddrBit),
				  CLKA => clk,
				  CLKB => clk,
				  DIA => memAWrite(31 downto 16),
				  DIB => memBWrite(31 downto 16),
				  DIPA => "00",
				  DIPB => "00",
				  ENA => '1',
				  ENB => '1',
				  SSRA => '0',
				  SSRB => '0',
				  WEA => memAWriteEnable,
				  WEB => memBWriteEnable);



	RAMB16_S18_S18_inst0: RAMB16_S18_S18
		generic map (
INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => x"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => x"0000000000000000000000000000000000000000000000000000000000000000")
		port map (DOA => memARead(15 downto 0),
				  DOB => memBRead(15 downto 0),
				  DOPA => open,
				  DOPB => open,
				  ADDRA => memAAddr(addrBitBRAM downto minAddrBit),
				  ADDRB => memBAddr(addrBitBRAM downto minAddrBit),
				  CLKA => clk,
				  CLKB => clk,
				  DIA => memAWrite(15 downto 0),
				  DIB => memBWrite(15 downto 0),
				  DIPA => "00",
				  DIPB => "00",
				  ENA => '1',
				  ENB => '1',
				  SSRA => '0',
				  SSRB => '0',
				  WEA => memAWriteEnable,
				  WEB => memBWriteEnable);
end behave_dualport_ram1;
